// Multiplexer testbench
`timescale 1 ns / 1 ps
`include "multiplexer.v"

module testMultiplexer ();
  reg address0, address1;
  reg in0, in1, in2, in3;
  wire out;

  // behavioralMultiplexer multiplexer (out, address0, address1, in0, in1, in2, in3);
  structuralMultiplexer multiplexer (out, address0, address1, in0, in1, in2, in3);

  initial begin
    $display("A0 A1 In0 In1 In2 In3 | Out | Expected Output");
    address0=0;address1=0;in0=1;in1=0;in2=0;in3=0; #1000
    $display("%b  %b   %b   %b   %b   %b  |  %b  | In0", address0, address1, in0, in1, in2, in3, out);
    address0=1;address1=0;in0=0;in1=1;in2=0;in3=0; #1000
    $display("%b  %b   %b   %b   %b   %b  |  %b  | In1", address0, address1, in0, in1, in2, in3, out);
    address0=0;address1=1;in0=0;in1=0;in2=1;in3=0; #1000
    $display("%b  %b   %b   %b   %b   %b  |  %b  | In2", address0, address1, in0, in1, in2, in3, out);
    address0=1;address1=1;in0=0;in1=0;in2=0;in3=1; #1000
    $display("%b  %b   %b   %b   %b   %b  |  %b  | In3", address0, address1, in0, in1, in2, in3, out);
    address0=0;address1=0;in0=0;in1=1;in2=1;in3=1; #1000
    $display("%b  %b   %b   %b   %b   %b  |  %b  | In0", address0, address1, in0, in1, in2, in3, out);
    address0=1;address1=0;in0=1;in1=0;in2=1;in3=1; #1000
    $display("%b  %b   %b   %b   %b   %b  |  %b  | In1", address0, address1, in0, in1, in2, in3, out);
    address0=0;address1=1;in0=1;in1=1;in2=0;in3=1; #1000
    $display("%b  %b   %b   %b   %b   %b  |  %b  | In2", address0, address1, in0, in1, in2, in3, out);
    address0=1;address1=1;in0=1;in1=1;in2=1;in3=0; #1000
    $display("%b  %b   %b   %b   %b   %b  |  %b  | In3", address0, address1, in0, in1, in2, in3, out);
  end
endmodule
